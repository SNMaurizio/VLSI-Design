magic
tech sky130A
magscale 1 2
timestamp 1648854593
<< nwell >>
rect 606 519 636 599
rect 1715 477 2293 507
rect 2425 -938 2435 -438
<< poly >>
rect 3141 653 3171 743
rect 3141 623 3264 653
rect 499 477 798 507
rect 589 -93 619 477
rect 887 287 917 543
rect 1045 503 1309 533
rect 1715 477 2293 507
rect 1805 -68 1835 302
rect 2417 -21 2447 305
rect 589 -123 713 -93
rect 1644 -98 1835 -68
rect 2387 -51 2447 -21
rect 3020 -33 3050 326
rect 3234 196 3264 623
rect 2387 -202 2417 -51
rect 3020 -63 3098 -33
rect 575 -497 605 -227
rect 2387 -232 2525 -202
rect 3068 -219 3098 -63
rect 3068 -249 3226 -219
rect 1107 -383 1275 -353
rect 2034 -489 2064 -290
rect 3044 -642 3074 -442
<< locali >>
rect 542 894 670 934
rect 1150 894 1278 934
rect 1758 894 1886 934
rect 2974 894 3098 934
rect 30 2 86 46
rect 566 2 646 46
rect 1174 2 1254 46
rect 2998 2 3074 46
rect 542 -886 670 -846
rect 1150 -886 1278 -846
rect 2366 -886 2494 -846
rect 2974 -886 3098 -846
<< metal1 >>
rect 4 696 105 752
rect 3122 744 3186 931
rect 284 481 428 511
rect 869 494 1525 524
rect 398 396 428 481
rect 398 366 1522 396
rect 2565 385 3084 415
rect 285 280 932 310
rect 589 -236 619 280
rect 1197 -184 1227 366
rect 1266 279 1853 309
rect 2581 106 2611 385
rect 1804 76 2611 106
rect 3020 156 3262 186
rect 1052 -214 1228 -184
rect 870 -307 1007 -306
rect 442 -336 1007 -307
rect 442 -337 897 -336
rect 977 -385 1007 -336
rect 1052 -385 1082 -214
rect 1643 -341 1673 -68
rect 1805 -288 1835 76
rect 2039 -277 2743 -247
rect 977 -414 1409 -385
rect 977 -415 2753 -414
rect 1379 -444 2753 -415
rect 904 -445 1351 -444
rect 162 -474 1351 -445
rect 3020 -461 3050 156
rect 3458 -150 3602 -94
rect 162 -475 904 -474
rect 1321 -488 1351 -474
rect 3181 -483 3502 -453
rect 1321 -518 2071 -488
rect 3181 -519 3211 -483
rect 2947 -549 3211 -519
rect 3030 -842 3087 -609
rect 3030 -890 3122 -842
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1648818724
transform 1 0 3040 0 1 -14
box -4 14 604 1000
use Inversor  Inversor_0 ~/icdesign/mag/Inversor
timestamp 1648821604
transform 1 0 608 0 1 2
box 0 -2 608 984
use Inversor  Inversor_1
timestamp 1648821604
transform 1 0 0 0 -1 46
box 0 -2 608 984
use Inversor  Inversor_2
timestamp 1648821604
transform 1 0 3036 0 -1 46
box 0 -2 608 984
use NOR  NOR_0 ~/icdesign/mag/NOR
timestamp 1648848246
transform -1 0 2467 0 -1 46
box 39 -2 1255 984
use NOR  NOR_1
timestamp 1648848246
transform 1 0 1785 0 1 2
box 39 -2 1255 984
use TGate  TGate_0 ~/icdesign/mag/TGate
timestamp 1648821211
transform 1 0 0 0 1 2
box 0 -2 608 984
use TGate  TGate_1
timestamp 1648821211
transform 1 0 608 0 -1 46
box 0 -2 608 984
use TGate  TGate_2
timestamp 1648821211
transform 1 0 1216 0 1 2
box 0 -2 608 984
use TGate  TGate_3
timestamp 1648821211
transform 1 0 2432 0 -1 46
box 0 -2 608 984
use via  via_0 ~/icdesign/mag/Via
timestamp 1647641870
transform 1 0 3407 0 1 -664
box 31 179 97 245
use via  via_1
timestamp 1647641870
transform 1 0 2995 0 1 -849
box 31 179 97 245
use via  via_2
timestamp 1647641870
transform 1 0 1756 0 1 68
box 31 179 97 245
use via  via_3
timestamp 1647641870
transform 1 0 1228 0 1 70
box 31 179 97 245
use via  via_4
timestamp 1647641870
transform 1 0 1757 0 1 -469
box 31 179 97 245
use via  via_5
timestamp 1647641870
transform 1 0 2531 0 1 174
box 31 179 97 245
use via  via_6
timestamp 1647641870
transform 1 0 3034 0 1 193
box 31 179 97 245
use via  via_7
timestamp 1647641870
transform 1 0 350 0 1 -549
box 31 179 97 245
use via  via_8
timestamp 1647641870
transform 1 0 834 0 1 -546
box 31 179 97 245
use via  via_9
timestamp 1647641870
transform 1 0 835 0 1 -659
box 31 179 97 245
use via  via_10
timestamp 1647641870
transform 1 0 129 0 1 -688
box 31 179 97 245
use via  via_11
timestamp 1647641870
transform 1 0 2001 0 1 -718
box 31 179 97 245
use via  via_12
timestamp 1647641870
transform 1 0 838 0 1 96
box 31 179 97 245
use via  via_13
timestamp 1647641870
transform 1 0 2659 0 1 -659
box 31 179 97 245
use via  via_14
timestamp 1647641870
transform 1 0 2658 0 1 -473
box 31 179 97 245
use via  via_15
timestamp 1647641870
transform 1 0 2000 0 1 -473
box 31 179 97 245
use via  via_16
timestamp 1647641870
transform 1 0 1430 0 1 156
box 31 179 97 245
use via  via_17
timestamp 1647641870
transform 1 0 1429 0 1 290
box 31 179 97 245
use via  via_18
timestamp 1647641870
transform 1 0 250 0 1 98
box 31 179 97 245
use via  via_19
timestamp 1647641870
transform 1 0 249 0 1 284
box 31 179 97 245
use via  via_20
timestamp 1647641870
transform 1 0 838 0 1 313
box 31 179 97 245
use via  via_21
timestamp 1647641870
transform 1 0 526 0 1 -690
box 31 179 97 245
use via  via_22
timestamp 1647641870
transform 1 0 526 0 1 -457
box 31 179 97 245
use via  via_23
timestamp 1647641870
transform 1 0 1597 0 1 -298
box 31 179 97 245
use via  via_24
timestamp 1647641870
transform 1 0 1594 0 1 -550
box 31 179 97 245
use via  via_25
timestamp 1647641870
transform 1 0 2984 0 1 -652
box 31 179 97 245
use via  via_26
timestamp 1647641870
transform 1 0 3185 0 1 -41
box 31 179 97 245
use via  via_27
timestamp 1647641870
transform 1 0 3091 0 1 557
box 31 179 97 245
<< labels >>
rlabel poly 3020 -63 3050 326 1 Q
rlabel space 3457 -150 3602 -94 1 Qb
rlabel space 176 -493 210 -459 1 clk
rlabel space 162 -475 931 -445 1 clk
rlabel metal1 4 696 105 752 1 D
rlabel space 2564 385 3084 415 1 clr
<< end >>
