magic
tech sky130A
magscale 1 2
timestamp 1648670410
<< nwell >>
rect 604 484 666 984
<< poly >>
rect 439 303 469 641
rect 794 386 824 622
rect 794 351 1110 386
rect 439 273 1022 303
rect 1080 267 1110 351
rect 1192 331 1222 561
<< metal1 >>
rect 95 677 140 928
rect 510 927 748 936
rect 193 641 237 815
rect 287 676 332 927
rect 479 888 748 927
rect 384 641 428 816
rect 479 676 524 888
rect 609 830 1169 860
rect 609 641 639 830
rect 740 657 781 830
rect 193 611 639 641
rect 836 622 878 795
rect 932 657 973 830
rect 1029 622 1069 798
rect 1125 659 1169 830
rect 836 592 1236 622
rect 1029 276 1234 332
rect 588 0 682 46
rect 943 8 983 243
rect 1029 101 1074 276
rect 1119 7 1159 242
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1647017803
transform 1 0 4 0 1 -16
box -4 16 604 1000
use 5umcell_template  5umcell_template_1
timestamp 1647017803
transform 1 0 666 0 1 -16
box -4 16 604 1000
use pfet_w075_4f  pfet_w075_4f_0 ~/icdesign/mag/PFET_W075_4f
timestamp 1647552966
transform 1 0 53 0 1 570
box 0 0 514 350
use pfet_w075_4f  pfet_w075_4f_1
timestamp 1647552966
transform 1 0 696 0 1 551
box 0 0 514 350
use sky130_fd_pr__nfet_01v8_SJ5Z6H  sky130_fd_pr__nfet_01v8_SJ5Z6H_0
timestamp 1648504841
transform 1 0 1007 0 1 173
box -73 -101 73 101
use sky130_fd_pr__nfet_01v8_SJ5Z6H  sky130_fd_pr__nfet_01v8_SJ5Z6H_1
timestamp 1648504841
transform 1 0 1095 0 1 173
box -73 -101 73 101
use via  via_0 ~/icdesign/mag/Via
timestamp 1647641870
transform 1 0 1141 0 1 376
box 31 179 97 245
use via  via_1
timestamp 1647641870
transform 1 0 1141 0 1 93
box 31 179 97 245
<< labels >>
rlabel space 98 894 498 930 1 Vdd
rlabel space 32 6 576 40 1 Vss
rlabel space 439 273 469 670 1 A
rlabel space 794 351 824 651 1 B
rlabel space 1192 322 1222 571 1 OUT
<< end >>
