magic
tech sky130A
magscale 1 2
timestamp 1647559469
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1647017803
transform 1 0 4 0 1 -16
box -4 16 604 1000
use nfet_w075_2f  nfet_w075_2f_0 ~/icdesign/mag/NFET_W075_2F
timestamp 1647552215
transform 1 0 -1145 0 1 -54
box 0 32 250 264
use nfet_w075_2f  nfet_w075_2f_1
timestamp 1647552215
transform 1 0 -620 0 1 -51
box 0 32 250 264
use pfet_w075_2f  pfet_w075_2f_0 ~/icdesign/mag/PFET_W075_2F
timestamp 1647552722
transform 1 0 -574 0 1 565
box 0 0 322 350
use pfet_w075_2f  pfet_w075_2f_1
timestamp 1647552722
transform 1 0 -1227 0 1 565
box 0 0 322 350
<< end >>
