* NGSPICE file created from Inversor.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_NDWVGB a_15_n75# a_n15_n101# a_n73_n75# VSUBS
X0 a_15_n75# a_n15_n101# a_n73_n75# VSUBS sky130_fd_pr__nfet_01v8 ad=2.175e+11p pd=2.08e+06u as=2.175e+11p ps=2.08e+06u w=750000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_52C9FB w_n161_n175# a_n63_n106# a_n33_n75# a_63_n75#
+ a_n125_n75#
X0 a_n33_n75# a_n63_n106# a_n125_n75# w_n161_n175# sky130_fd_pr__pfet_01v8 ad=2.475e+11p pd=2.16e+06u as=2.325e+11p ps=2.12e+06u w=750000u l=150000u
X1 a_63_n75# a_n63_n106# a_n33_n75# w_n161_n175# sky130_fd_pr__pfet_01v8 ad=2.325e+11p pd=2.12e+06u as=0p ps=0u w=750000u l=150000u
.ends

.subckt pfet_w075_2f sky130_fd_pr__pfet_01v8_52C9FB_0/a_n33_n75# sky130_fd_pr__pfet_01v8_52C9FB_0/a_63_n75#
+ sky130_fd_pr__pfet_01v8_52C9FB_0/a_n125_n75# sky130_fd_pr__pfet_01v8_52C9FB_0/w_n161_n175#
+ sky130_fd_pr__pfet_01v8_52C9FB_0/a_n63_n106#
Xsky130_fd_pr__pfet_01v8_52C9FB_0 sky130_fd_pr__pfet_01v8_52C9FB_0/w_n161_n175# sky130_fd_pr__pfet_01v8_52C9FB_0/a_n63_n106#
+ sky130_fd_pr__pfet_01v8_52C9FB_0/a_n33_n75# sky130_fd_pr__pfet_01v8_52C9FB_0/a_63_n75#
+ sky130_fd_pr__pfet_01v8_52C9FB_0/a_n125_n75# sky130_fd_pr__pfet_01v8_52C9FB
.ends


* Top level circuit Inversor

Xsky130_fd_pr__nfet_01v8_NDWVGB_0 m1_200_106# a_160_274# VSUBS VSUBS sky130_fd_pr__nfet_01v8_NDWVGB
Xpfet_w075_2f_0 m1_200_106# m1_299_677# m1_299_677# m1_299_677# a_160_274# pfet_w075_2f
.end

