magic
tech sky130A
magscale 1 2
timestamp 1648848246
<< poly >>
rect 478 303 508 641
rect 794 386 824 622
rect 794 351 1110 386
rect 478 273 1022 303
rect 1080 267 1110 351
rect 1192 331 1222 561
<< locali >>
rect 581 892 709 932
rect 605 0 685 44
<< metal1 >>
rect 134 677 179 928
rect 232 641 276 815
rect 326 676 371 927
rect 423 641 467 816
rect 518 670 563 936
rect 632 830 1169 860
rect 632 641 662 830
rect 740 657 781 830
rect 232 611 662 641
rect 836 622 878 795
rect 932 657 973 830
rect 1029 622 1069 798
rect 1125 659 1169 830
rect 836 592 1236 622
rect 1029 295 1234 351
rect 943 8 983 243
rect 1029 101 1074 295
rect 1119 7 1159 242
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1648818724
transform 1 0 43 0 1 -16
box -4 14 604 1000
use 5umcell_template  5umcell_template_1
timestamp 1648818724
transform 1 0 651 0 1 -16
box -4 14 604 1000
use pfet_w075_4f  pfet_w075_4f_0 ~/icdesign/mag/PFET_W075_4f
timestamp 1647552966
transform 1 0 92 0 1 570
box 0 0 514 350
use pfet_w075_4f  pfet_w075_4f_1
timestamp 1647552966
transform 1 0 696 0 1 551
box 0 0 514 350
use sky130_fd_pr__nfet_01v8_SJ5Z6H  sky130_fd_pr__nfet_01v8_SJ5Z6H_2
timestamp 1648817418
transform 1 0 1007 0 1 173
box -73 -101 73 101
use sky130_fd_pr__nfet_01v8_SJ5Z6H  sky130_fd_pr__nfet_01v8_SJ5Z6H_3
timestamp 1648817418
transform 1 0 1095 0 1 173
box -73 -101 73 101
use via  via_0 ~/icdesign/mag/Via
timestamp 1647641870
transform 1 0 1141 0 1 376
box 31 179 97 245
use via  via_1
timestamp 1647641870
transform 1 0 1141 0 1 112
box 31 179 97 245
<< labels >>
rlabel space 794 351 824 651 1 B
rlabel space 478 273 508 670 1 A
rlabel space 137 894 537 930 1 Vdd
rlabel space 747 4 1147 40 1 Vss
rlabel space 1192 331 1222 571 1 OUT
<< end >>
