* NGSPICE file created from NAND.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_XUMWGH a_n33_n75# a_63_n75# a_n125_n75# a_n63_n131#
+ VSUBS
X0 a_63_n75# a_n63_n131# a_n33_n75# VSUBS sky130_fd_pr__nfet_01v8 ad=2.325e+11p pd=2.12e+06u as=2.475e+11p ps=2.16e+06u w=750000u l=150000u
X1 a_n33_n75# a_n63_n131# a_n125_n75# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.325e+11p ps=2.12e+06u w=750000u l=150000u
.ends

.subckt nfet_w075_2f sky130_fd_pr__nfet_01v8_XUMWGH_0/a_n125_n75# sky130_fd_pr__nfet_01v8_XUMWGH_0/a_n63_n131#
+ sky130_fd_pr__nfet_01v8_XUMWGH_0/a_n33_n75# sky130_fd_pr__nfet_01v8_XUMWGH_0/a_63_n75#
Xsky130_fd_pr__nfet_01v8_XUMWGH_0 sky130_fd_pr__nfet_01v8_XUMWGH_0/a_n33_n75# sky130_fd_pr__nfet_01v8_XUMWGH_0/a_63_n75#
+ sky130_fd_pr__nfet_01v8_XUMWGH_0/a_n125_n75# sky130_fd_pr__nfet_01v8_XUMWGH_0/a_n63_n131#
+ VSUBS sky130_fd_pr__nfet_01v8_XUMWGH
.ends

.subckt sky130_fd_pr__pfet_01v8_52C9FB w_n161_n175# a_n63_n106# a_n33_n75# a_63_n75#
+ a_n125_n75#
X0 a_n33_n75# a_n63_n106# a_n125_n75# w_n161_n175# sky130_fd_pr__pfet_01v8 ad=2.475e+11p pd=2.16e+06u as=2.325e+11p ps=2.12e+06u w=750000u l=150000u
X1 a_63_n75# a_n63_n106# a_n33_n75# w_n161_n175# sky130_fd_pr__pfet_01v8 ad=2.325e+11p pd=2.12e+06u as=0p ps=0u w=750000u l=150000u
.ends

.subckt pfet_w075_2f sky130_fd_pr__pfet_01v8_52C9FB_0/a_n33_n75# sky130_fd_pr__pfet_01v8_52C9FB_0/a_63_n75#
+ sky130_fd_pr__pfet_01v8_52C9FB_0/a_n125_n75# sky130_fd_pr__pfet_01v8_52C9FB_0/w_n161_n175#
+ sky130_fd_pr__pfet_01v8_52C9FB_0/a_n63_n106#
Xsky130_fd_pr__pfet_01v8_52C9FB_0 sky130_fd_pr__pfet_01v8_52C9FB_0/w_n161_n175# sky130_fd_pr__pfet_01v8_52C9FB_0/a_n63_n106#
+ sky130_fd_pr__pfet_01v8_52C9FB_0/a_n33_n75# sky130_fd_pr__pfet_01v8_52C9FB_0/a_63_n75#
+ sky130_fd_pr__pfet_01v8_52C9FB_0/a_n125_n75# sky130_fd_pr__pfet_01v8_52C9FB
.ends


* Top level circuit NAND

Xnfet_w075_2f_0 m1_32_136# a_86_283# VSUBS m1_32_136# nfet_w075_2f
Xnfet_w075_2f_1 OUT a_392_299# m1_32_136# OUT nfet_w075_2f
Xpfet_w075_2f_0 OUT m1_87_677# m1_87_677# m1_87_677# a_86_283# pfet_w075_2f
Xpfet_w075_2f_1 OUT m1_87_677# m1_87_677# m1_87_677# a_392_299# pfet_w075_2f
.end

