magic
tech sky130A
timestamp 1647004767
<< nwell >>
rect 0 250 300 500
<< psubdiff >>
rect -2 10 10 30
rect 290 10 302 30
<< nsubdiff >>
rect 25 473 273 474
rect 25 455 47 473
rect 247 455 273 473
rect 25 454 273 455
<< psubdiffcont >>
rect 10 10 290 30
<< nsubdiffcont >>
rect 47 455 247 473
<< locali >>
rect 29 473 269 474
rect 29 455 47 473
rect 247 455 269 473
rect 29 454 269 455
rect 2 10 10 30
rect 290 10 298 30
<< end >>
