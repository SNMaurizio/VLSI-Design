magic
tech sky130A
magscale 1 2
timestamp 1647646778
<< nwell >>
rect 67 533 132 1033
<< poly >>
rect -461 352 -414 690
rect -153 352 -106 690
<< metal1 >>
rect -504 981 36 984
rect -504 938 226 981
rect -504 936 36 938
rect -504 724 -456 936
rect -411 688 -361 865
rect -320 720 -272 936
rect -204 724 -156 936
rect -106 688 -56 865
rect -12 722 36 936
rect -411 658 61 688
rect -1 493 50 658
rect -1 445 286 493
rect -518 388 -52 397
rect -519 369 -50 388
rect -519 186 -468 369
rect -424 65 -373 324
rect -328 183 -277 369
rect -192 150 -145 322
rect -101 186 -50 369
rect -1 182 50 445
rect 0 150 47 182
rect -192 122 47 150
rect 48 50 163 93
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1647017803
transform 1 0 -533 0 1 32
box -4 16 604 1000
use Inversor  Inversor_0 ~/icdesign/mag/Inversor
timestamp 1647642706
transform 1 0 128 0 1 49
box 0 0 608 984
use nfet_w075_2f  nfet_w075_2f_0 ~/icdesign/mag/NFET_W075_2F
timestamp 1647552215
transform 1 0 -523 0 1 90
box 0 32 250 264
use nfet_w075_2f  nfet_w075_2f_1
timestamp 1647552215
transform 1 0 -198 0 1 90
box 0 32 250 264
use pfet_w075_2f  pfet_w075_2f_0 ~/icdesign/mag/PFET_W075_2F
timestamp 1647552722
transform 1 0 -245 0 1 618
box 0 0 322 350
use pfet_w075_2f  pfet_w075_2f_1
timestamp 1647552722
transform 1 0 -549 0 1 618
box 0 0 322 350
use via  via_0 ~/icdesign/mag/Via
timestamp 1647641870
transform 1 0 192 0 1 259
box 31 179 97 245
<< labels >>
rlabel poly -461 352 -414 690 1 B
rlabel poly -153 352 -106 690 1 A
rlabel space 328 155 372 869 1 OUT
<< end >>
