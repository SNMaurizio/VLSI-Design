* NGSPICE file created from /home/designer/icdesign/mag/inv/Inversor.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_PDE3P4 a_n33_36# a_15_n76# a_n73_n76# VSUBS
X0 a_15_n76# a_n33_36# a_n73_n76# VSUBS sky130_fd_pr__nfet_01v8 ad=1.305e+11p pd=1.48e+06u as=1.305e+11p ps=1.48e+06u w=450000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_A9BS5R a_n73_n9# a_15_n9# a_n33_n106# w_n109_n109#
X0 a_15_n9# a_n33_n106# a_n73_n9# w_n109_n109# sky130_fd_pr__pfet_01v8 ad=1.305e+11p pd=1.48e+06u as=1.305e+11p ps=1.48e+06u w=450000u l=150000u
.ends


* Top level circuit /home/designer/icdesign/mag/inv/Inversor

Xsky130_fd_pr__nfet_01v8_PDE3P4_0 IN OUT sky130_fd_pr__pfet_01v8_A9BS5R_0/VSUBS sky130_fd_pr__pfet_01v8_A9BS5R_0/VSUBS
+ sky130_fd_pr__nfet_01v8_PDE3P4
Xsky130_fd_pr__pfet_01v8_A9BS5R_0 Vdd OUT IN Vdd sky130_fd_pr__pfet_01v8_A9BS5R
.end

