magic
tech sky130A
magscale 1 2
timestamp 1649112742
<< nwell >>
rect 4238 972 4264 1437
rect 4243 -2811 4261 -2311
<< poly >>
rect 3487 147 3768 188
rect 3842 157 4384 187
rect 3490 -138 4035 -108
<< metal1 >>
rect 3731 2708 3782 2815
rect 3280 2253 4612 2306
rect 3401 2179 3516 2221
rect 3737 2040 3789 2253
rect 4377 2179 4492 2221
rect 3727 1988 3737 2040
rect 3789 1988 3799 2040
rect 3671 1875 3751 1923
rect 4078 1877 4129 1984
rect 3727 1771 3737 1823
rect 3789 1771 3799 1823
rect 90 1373 100 1425
rect 152 1373 162 1425
rect 3737 1148 3789 1771
rect 7733 1373 7743 1425
rect 7795 1373 7805 1425
rect 3727 1096 3737 1148
rect 3789 1096 3799 1148
rect 6031 937 6041 989
rect 6093 937 6103 989
rect 3727 791 3737 843
rect 3789 831 3799 843
rect 3789 801 4154 831
rect 3789 791 3799 801
rect 3553 320 3594 434
rect 3714 306 3724 358
rect 3776 306 3786 358
rect 3728 145 3758 306
rect 3819 137 3829 189
rect 3881 137 3891 189
rect 4124 157 4154 801
rect 4307 309 4317 361
rect 4369 309 4379 361
rect 4104 105 4114 157
rect 4166 105 4176 157
rect 3671 1 3751 49
rect 4104 -80 4114 -28
rect 4166 -80 4176 -28
rect 3989 -147 3999 -95
rect 4051 -147 4061 -95
rect 3533 -312 3543 -260
rect 3595 -312 3605 -260
rect 4133 -751 4163 -80
rect 4292 -310 4302 -258
rect 4354 -310 4364 -258
rect 4110 -803 4120 -751
rect 4172 -803 4182 -751
rect 6031 -938 6041 -886
rect 6093 -938 6103 -886
rect 4110 -1066 4120 -1014
rect 4172 -1066 4182 -1014
rect 89 -1375 99 -1323
rect 151 -1375 161 -1323
rect 104 -1468 134 -1375
rect 4136 -1672 4166 -1066
rect 7736 -1376 7746 -1324
rect 7798 -1376 7808 -1324
rect 4111 -1724 4121 -1672
rect 4173 -1724 4183 -1672
rect 3645 -1874 3765 -1825
rect 4144 -1875 4264 -1826
rect 4111 -1958 4121 -1906
rect 4173 -1958 4183 -1906
rect 3402 -2171 3521 -2129
rect 4121 -2203 4173 -1958
rect 4373 -2171 4492 -2129
rect 3281 -2256 4620 -2203
<< via1 >>
rect 3737 1988 3789 2040
rect 3737 1771 3789 1823
rect 100 1373 152 1425
rect 7743 1373 7795 1425
rect 3737 1096 3789 1148
rect 6041 937 6093 989
rect 3737 791 3789 843
rect 3724 306 3776 358
rect 3829 137 3881 189
rect 4317 309 4369 361
rect 4114 105 4166 157
rect 4114 -80 4166 -28
rect 3999 -147 4051 -95
rect 3543 -312 3595 -260
rect 4302 -310 4354 -258
rect 4120 -803 4172 -751
rect 6041 -938 6093 -886
rect 4120 -1066 4172 -1014
rect 99 -1375 151 -1323
rect 7746 -1376 7798 -1324
rect 4121 -1724 4173 -1672
rect 4121 -1958 4173 -1906
<< metal2 >>
rect 3737 2040 3789 2050
rect 3737 1978 3789 1988
rect 3737 1833 3788 1978
rect 3737 1823 3789 1833
rect 3737 1761 3789 1771
rect 100 1425 152 1435
rect 7743 1425 7795 1435
rect 10 1373 100 1425
rect 152 1373 7743 1425
rect 7795 1373 7888 1425
rect 10 -1324 40 1373
rect 100 1363 152 1373
rect 7743 1363 7795 1373
rect 3737 1148 3789 1158
rect 3737 843 3789 1096
rect 3737 781 3789 791
rect 6041 989 6093 999
rect 3724 358 3776 368
rect 4317 361 4369 371
rect 3776 318 4317 348
rect 3724 296 3776 306
rect 4317 299 4369 309
rect 3829 189 3881 199
rect 3829 127 3881 137
rect 4114 157 4166 167
rect 3543 -260 3595 -250
rect 3845 -269 3874 127
rect 4114 -28 4166 105
rect 3999 -95 4051 -85
rect 4114 -90 4166 -80
rect 3999 -157 4051 -147
rect 3595 -298 3874 -269
rect 4013 -272 4041 -157
rect 4302 -258 4354 -248
rect 4013 -300 4302 -272
rect 3543 -322 3595 -312
rect 4302 -320 4354 -310
rect 4120 -751 4172 -741
rect 4120 -1014 4172 -803
rect 6041 -886 6093 937
rect 6041 -948 6093 -938
rect 4120 -1076 4172 -1066
rect 99 -1323 151 -1313
rect 10 -1375 99 -1324
rect 10 -1376 151 -1375
rect 99 -1385 151 -1376
rect 7746 -1324 7798 -1314
rect 7858 -1324 7888 1373
rect 7798 -1376 7888 -1324
rect 7746 -1386 7798 -1376
rect 4121 -1672 4173 -1662
rect 4121 -1906 4173 -1724
rect 4121 -1968 4173 -1958
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1648818724
transform 1 0 3648 0 1 1861
box -4 14 604 1000
use 5umcell_template  5umcell_template_1
timestamp 1648818724
transform -1 0 4244 0 -1 1937
box -4 14 604 1000
use 5umcell_template  5umcell_template_2
timestamp 1648818724
transform 1 0 3652 0 1 -13
box -4 14 604 1000
use 5umcell_template  5umcell_template_3
timestamp 1648818724
transform -1 0 4248 0 -1 63
box -4 14 604 1000
use 5umcell_template  5umcell_template_4
timestamp 1648818724
transform 1 0 3648 0 1 -1887
box -4 14 604 1000
use 5umcell_template  5umcell_template_5
timestamp 1648818724
transform -1 0 4244 0 -1 -1811
box -4 14 604 1000
use contador_1bit  contador_1bit_0 ~/icdesign/mag/Contador1bit
timestamp 1649101816
transform 1 0 1901 0 1 -481
box -1901 481 1784 3342
use contador_1bit  contador_1bit_1
timestamp 1649101816
transform -1 0 5995 0 1 -481
box -1901 481 1784 3342
use contador_1bit  contador_1bit_2
timestamp 1649101816
transform 1 0 1901 0 -1 531
box -1901 481 1784 3342
use contador_1bit  contador_1bit_3
timestamp 1649101816
transform -1 0 5995 0 -1 531
box -1901 481 1784 3342
use via  via_0 ~/icdesign/mag/Via
timestamp 1647641870
transform 1 0 3680 0 1 -47
box 31 179 97 245
use via  via_1
timestamp 1647641870
transform 1 0 3790 0 1 -49
box 31 179 97 245
use via  via_2
timestamp 1647641870
transform 1 0 3962 0 1 -335
box 31 179 97 245
<< labels >>
rlabel metal1 3553 320 3594 434 1 CE
rlabel metal1 3731 2708 3782 2815 1 VDD
rlabel metal1 4078 1877 4129 1984 1 VSS
rlabel metal1 3401 2179 3516 2221 1 D0
rlabel metal1 4377 2179 4492 2221 1 D1
rlabel metal1 3402 -2171 3521 -2129 1 D2
rlabel metal1 4373 -2171 4492 -2129 1 D3
rlabel metal1 3737 2040 3789 2306 1 CLR
rlabel metal1 104 -1468 134 -1344 1 CLK
<< end >>
