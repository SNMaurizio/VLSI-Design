magic
tech sky130A
magscale 1 2
timestamp 1648821604
<< poly >>
rect 160 851 286 881
rect 160 274 190 639
rect 437 201 467 576
<< metal1 >>
rect 107 674 147 924
rect 203 629 243 813
rect 299 677 339 927
rect 203 581 474 629
rect 112 6 150 241
rect 200 194 239 247
rect 196 141 479 194
rect 200 101 239 141
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1648818724
transform 1 0 4 0 1 -16
box -4 14 604 1000
use pfet_w075_2f  pfet_w075_2f_0 ~/icdesign/mag/PFET_W075_2F
timestamp 1648666716
transform 1 0 62 0 1 570
box 0 0 322 350
use sky130_fd_pr__nfet_01v8_NDWVGB  sky130_fd_pr__nfet_01v8_NDWVGB_0
timestamp 1647553962
transform 1 0 175 0 1 175
box -73 -101 73 101
use via  via_0 ~/icdesign/mag/Via
timestamp 1647641870
transform 1 0 388 0 1 394
box 31 179 97 245
use via  via_1
timestamp 1647641870
transform 1 0 388 0 1 -43
box 31 179 97 245
<< labels >>
rlabel space 160 248 190 670 1 IN
rlabel space 98 894 498 930 1 Vdd
rlabel space 437 186 467 589 1 OUT
rlabel space 100 4 500 40 1 Vss
<< end >>
