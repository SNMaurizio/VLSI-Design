** sch_path: /home/designer/icdesign/sch//NMOS/Ej1.sch
**.subckt Ej1
XM1 d g GND GND sky130_fd_pr__nfet_01v8 L=3 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
VGS g GND DC{vgs}
VDS d GND DC{vds}
**** begin user architecture code



* Parameters
.param vds = 1.8
.param vgs = 0.9
.options TEMPS = 27.0

* Models
.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib TT

* Data to save
.save all  @M.XM1.msky130_fd_pr__nfet_01v8[id]  @M.XM1.msky130_fd_pr__nfet_01v8[gm]  @M.XM1.msky130_fd_pr__nfet_01v8[vth]  @M.XM1.msky130_fd_pr__nfet_01v8[vds]  @M.XM1.msky130_fd_pr__nfet_01v8[vdsat]  @M.XM1.msky130_fd_pr__nfet_01v8[vgs]


* Simulation
.control
  dc VDS 0 1.8 0.01 VGS 0 1.8 0.3
  setplot dc1
  plot @M.XM1.msky130_fd_pr__nfet_01v8[id] ylabel Id xlabel Vds title 'Id vs Vds vs Vgs'
  set filetype = ascii
  write tp1_1_dc1.raw
.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
