** sch_path: /home/designer/icdesign/sch//And/tb_AND.sch
**.subckt tb_AND
V1 Vss GND DC{vss}
V2 Vdd Vss DC{vdd}
V3 INA Vss PULSE({vdd} {vss} 0 1p 1p {TClk/4} {TClk/2})DC 0 AC 0
V4 INB Vss PULSE({vdd} {vss} {TClk/8} 1p 1p {TClk/4} {TClk/2})DC 0 AC 0
x1 outAND Vdd INA INB Vss AND
**** begin user architecture code





* Circuit Parameters
.param vdd  = 1.8
.param vss  = 0.0
.param Tclk = 10n
.options TEMP = 65.0


* Include Models
.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib TT


* OP Parameters & Singals to save
.save all


*Simulations
.control
  tran 0.01u 100n
  setplot tran1
  plot v(INA)v(INB)+2 v(outAND)+4
.endc
.end


**** end user architecture code
**.ends

* expanding   symbol:  And/AND.sym # of pins=5
** sym_path: /home/designer/icdesign/sch//And/AND.sym
** sch_path: /home/designer/icdesign/sch//And/AND.sch
.subckt AND  OUT Vdd A B Vss
*.ipin Vss
*.ipin Vdd
*.ipin A
*.opin OUT
*.ipin B
x1 Vdd A B net1 Vss NAND
x2 Vdd net1 OUT Vss Inversor
.ends


* expanding   symbol:  NAND/NAND.sym # of pins=5
** sym_path: /home/designer/icdesign/sch//NAND/NAND.sym
** sch_path: /home/designer/icdesign/sch//NAND/NAND.sch
.subckt NAND  Vdd A B OUT Vss
*.ipin A
*.ipin B
*.ipin Vdd
*.ipin Vss
*.opin OUT
XM1 net1 B Vss Vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM2 OUT A net1 Vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM5 OUT B Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM4 OUT A Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  Inversor/Inversor.sym # of pins=4
** sym_path: /home/designer/icdesign/sch//Inversor/Inversor.sym
** sch_path: /home/designer/icdesign/sch//Inversor/Inversor.sch
.subckt Inversor  Vdd IN OUT Vss
*.ipin IN
*.ipin Vdd
*.ipin Vss
*.opin OUT
XM1 OUT IN Vss Vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends

.GLOBAL GND
.end
