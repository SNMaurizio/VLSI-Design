magic
tech sky130A
magscale 1 2
timestamp 1646770120
<< error_p >>
rect -29 -56 29 -50
rect -29 -90 -17 -56
rect -29 -96 29 -90
<< nwell >>
rect -109 -109 109 143
<< pmos >>
rect -15 -9 15 81
<< pdiff >>
rect -73 69 -15 81
rect -73 3 -61 69
rect -27 3 -15 69
rect -73 -9 -15 3
rect 15 69 73 81
rect 15 3 27 69
rect 61 3 73 69
rect 15 -9 73 3
<< pdiffc >>
rect -61 3 -27 69
rect 27 3 61 69
<< poly >>
rect -15 81 15 107
rect -15 -40 15 -9
rect -33 -56 33 -40
rect -33 -90 -17 -56
rect 17 -90 33 -56
rect -33 -106 33 -90
<< polycont >>
rect -17 -90 17 -56
<< locali >>
rect -61 69 -27 85
rect -61 -13 -27 3
rect 27 69 61 85
rect 27 -13 61 3
rect -33 -90 -17 -56
rect 17 -90 33 -56
<< viali >>
rect -61 3 -27 69
rect 27 3 61 69
rect -17 -90 17 -56
<< metal1 >>
rect -67 69 -21 81
rect -67 3 -61 69
rect -27 3 -21 69
rect -67 -9 -21 3
rect 21 69 67 81
rect 21 3 27 69
rect 61 3 67 69
rect 21 -9 67 3
rect -29 -56 29 -50
rect -29 -90 -17 -56
rect 17 -90 29 -56
rect -29 -96 29 -90
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.45 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
