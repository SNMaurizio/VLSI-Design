magic
tech sky130A
timestamp 1647017803
<< nwell >>
rect 0 250 300 500
<< psubdiff >>
rect -2 10 10 30
rect 290 10 302 30
<< nsubdiff >>
rect 25 473 273 474
rect 25 455 47 473
rect 247 455 273 473
rect 25 454 273 455
<< psubdiffcont >>
rect 10 10 290 30
<< nsubdiffcont >>
rect 47 455 247 473
<< locali >>
rect 29 473 269 474
rect 29 455 47 473
rect 247 455 269 473
rect 29 454 269 455
rect 2 10 10 30
rect 290 10 298 30
<< viali >>
rect 47 455 247 473
rect 14 11 286 28
<< metal1 >>
rect 41 473 253 476
rect 41 455 47 473
rect 247 455 253 473
rect 41 452 253 455
rect 8 28 292 31
rect 8 11 14 28
rect 286 11 292 28
rect 8 8 292 11
<< end >>
