magic
tech sky130A
magscale 1 2
timestamp 1648591444
<< nwell >>
rect -831 484 -768 984
rect -168 484 -105 984
rect 495 899 558 984
rect 495 484 558 549
<< poly >>
rect 905 382 935 513
<< metal1 >>
rect -927 888 -684 936
rect -264 888 -21 936
rect 94 621 133 795
rect 189 652 230 928
rect 401 888 640 936
rect 284 828 519 858
rect 284 621 328 828
rect 94 591 328 621
rect 382 563 425 795
rect 478 621 519 828
rect 573 654 614 888
rect 671 828 905 858
rect 671 621 714 828
rect 478 591 714 621
rect 764 563 807 791
rect 862 655 905 828
rect 382 533 950 563
rect 249 368 766 398
rect -40 310 193 340
rect -40 132 3 310
rect -849 0 -750 46
rect -186 0 -87 46
rect 54 9 97 282
rect 150 104 193 310
rect 249 138 289 368
rect 736 352 766 368
rect 475 310 708 340
rect 736 322 950 352
rect 345 104 385 282
rect 475 138 518 310
rect 150 74 385 104
rect 570 46 613 278
rect 665 104 708 310
rect 762 137 803 322
rect 860 104 900 275
rect 665 74 900 104
rect 479 9 613 46
rect 479 0 574 9
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1647017803
transform 1 0 -105 0 1 -16
box -4 16 604 1000
use 5umcell_template  5umcell_template_1
timestamp 1647017803
transform 1 0 558 0 1 -16
box -4 16 604 1000
use Inversor  Inversor_0 ~/icdesign/mag/Inversor
timestamp 1648588024
transform 1 0 -772 0 1 0
box 0 0 608 984
use Inversor  Inversor_1
timestamp 1648588024
transform 1 0 -1435 0 1 0
box 0 0 608 984
use pfet_w075_2f  pfet_w075_2f_0 ~/icdesign/mag/PFET_W075_2F
timestamp 1647552722
transform 1 0 49 0 1 549
box 0 0 322 350
use pfet_w075_2f  pfet_w075_2f_1
timestamp 1647552722
transform 1 0 241 0 1 549
box 0 0 322 350
use pfet_w075_2f  pfet_w075_2f_2
timestamp 1647552722
transform 1 0 433 0 1 549
box 0 0 322 350
use pfet_w075_2f  pfet_w075_2f_3
timestamp 1647552722
transform 1 0 625 0 1 549
box 0 0 322 350
use sky130_fd_pr__nfet_01v8_XE8V5F  sky130_fd_pr__nfet_01v8_XE8V5F_0
timestamp 1648583825
transform 1 0 76 0 1 207
box -125 -131 125 101
use sky130_fd_pr__nfet_01v8_XE8V5F  sky130_fd_pr__nfet_01v8_XE8V5F_1
timestamp 1648583825
transform 1 0 268 0 1 207
box -125 -131 125 101
use sky130_fd_pr__nfet_01v8_XE8V5F  sky130_fd_pr__nfet_01v8_XE8V5F_2
timestamp 1648583825
transform 1 0 783 0 1 207
box -125 -131 125 101
use sky130_fd_pr__nfet_01v8_XE8V5F  sky130_fd_pr__nfet_01v8_XE8V5F_3
timestamp 1648583825
transform 1 0 591 0 1 207
box -125 -131 125 101
use via  via_0 ~/icdesign/mag/Via
timestamp 1647641870
transform 1 0 213 0 1 1027
box 31 179 97 245
use via  via_1
timestamp 1647641870
transform 1 0 68 0 1 1023
box 31 179 97 245
use via  via_2
timestamp 1647641870
transform -1 0 984 0 -1 563
box 31 179 97 245
use via  via_3
timestamp 1647641870
transform 1 0 856 0 1 331
box 31 179 97 245
<< labels >>
rlabel space -85 4 475 44 1 Vss
rlabel space -11 894 389 930 1 Vdd
<< end >>
