magic
tech sky130A
magscale 1 2
timestamp 1647552722
<< nwell >>
rect -161 -175 161 175
<< pmos >>
rect -63 -75 -33 75
rect 33 -75 63 75
<< pdiff >>
rect -125 63 -63 75
rect -125 -63 -113 63
rect -79 -63 -63 63
rect -125 -75 -63 -63
rect -33 63 33 75
rect -33 -63 -17 63
rect 17 -63 33 63
rect -33 -75 33 -63
rect 63 63 125 75
rect 63 -63 79 63
rect 113 -63 125 63
rect 63 -75 125 -63
<< pdiffc >>
rect -113 -63 -79 63
rect -17 -63 17 63
rect 79 -63 113 63
<< poly >>
rect -63 106 63 136
rect -63 75 -33 106
rect 33 75 63 106
rect -63 -106 -33 -75
rect 33 -106 63 -75
<< locali >>
rect -113 63 -79 79
rect -113 -79 -79 -63
rect -17 63 17 79
rect -17 -79 17 -63
rect 79 63 113 79
rect 79 -79 113 -63
<< viali >>
rect -113 -63 -79 63
rect -17 -63 17 63
rect 79 -63 113 63
<< metal1 >>
rect -119 63 -73 75
rect -119 -63 -113 63
rect -79 -63 -73 63
rect -119 -75 -73 -63
rect -23 63 23 75
rect -23 -63 -17 63
rect 17 -63 23 63
rect -23 -75 23 -63
rect 73 63 119 75
rect 73 -63 79 63
rect 113 -63 119 63
rect 73 -75 119 -63
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.75 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
