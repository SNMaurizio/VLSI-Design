magic
tech sky130A
magscale 1 2
timestamp 1648483063
<< nwell >>
rect 67 533 132 1033
<< poly >>
rect -393 443 -363 718
rect -461 413 -363 443
rect -105 443 -75 690
rect -105 413 -10 443
rect -461 353 -431 413
rect -40 353 -10 413
<< metal1 >>
rect -456 936 -320 984
rect -272 941 -204 984
rect -272 936 -208 941
rect -156 936 235 984
rect -451 726 -401 936
rect -355 688 -307 867
rect -258 724 -208 936
rect -161 688 -113 867
rect -68 726 -18 936
rect -355 658 50 688
rect -1 493 50 658
rect -1 445 286 493
rect -519 369 -50 397
rect -519 186 -468 369
rect -424 65 -373 324
rect -328 183 -277 369
rect -192 150 -145 322
rect -101 186 -50 369
rect -1 182 50 445
rect 0 150 47 182
rect -192 122 47 150
rect 48 50 163 93
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1647017803
transform 1 0 -533 0 1 32
box -4 16 604 1000
use Inversor  Inversor_0 ~/icdesign/mag/Inversor
timestamp 1647647265
transform 1 0 128 0 1 49
box 0 0 608 984
use nfet_w075_2f  nfet_w075_2f_0 ~/icdesign/mag/NFET_W075_2F
timestamp 1647552215
transform 1 0 -523 0 1 90
box 0 32 250 264
use nfet_w075_2f  nfet_w075_2f_1
timestamp 1647552215
transform 1 0 -198 0 1 90
box 0 32 250 264
use pfet_w075_2f  pfet_w075_2f_0 ~/icdesign/mag/PFET_W075_2F
timestamp 1647552722
transform 1 0 -299 0 1 618
box 0 0 322 350
use pfet_w075_2f  pfet_w075_2f_1
timestamp 1647552722
transform 1 0 -491 0 1 618
box 0 0 322 350
use via  via_0 ~/icdesign/mag/Via
timestamp 1647641870
transform 1 0 192 0 1 259
box 31 179 97 245
<< labels >>
rlabel space 328 155 372 869 1 OUT
rlabel space -105 413 -75 718 1 A
rlabel poly -393 413 -363 718 1 B
<< end >>
