magic
tech sky130A
magscale 1 2
timestamp 1648496806
<< poly >>
rect 154 471 184 613
rect 155 274 185 416
<< metal1 >>
rect 100 822 336 859
rect 101 791 143 822
rect 101 102 145 791
rect 194 102 238 791
rect 292 648 334 822
use 5umcell_template  5umcell_template_0 ~/icdesign/mag/Plantilla
timestamp 1647017803
transform 1 0 4 0 1 -16
box -4 16 604 1000
use pfet_w075_2f  pfet_w075_2f_0 ~/icdesign/mag/PFET_W075_2F
timestamp 1647552722
transform 1 0 56 0 1 544
box 0 0 322 350
use sky130_fd_pr__nfet_01v8_SJ5Z6H  sky130_fd_pr__nfet_01v8_SJ5Z6H_0
timestamp 1647557214
transform 1 0 170 0 1 173
box -73 -101 73 101
<< labels >>
rlabel metal1 101 102 145 791 1 IN
rlabel metal1 194 102 238 791 1 OUT
rlabel space 154 471 184 644 1 Eb
rlabel space 155 248 185 416 1 E
rlabel space 98 894 498 930 1 Vdd
rlabel space 32 6 576 40 1 Vss
<< end >>
