magic
tech sky130A
magscale 1 2
timestamp 1648589124
<< nwell >>
rect 277 962 339 1462
<< metal1 >>
rect 185 1366 427 1414
rect 53 895 492 951
rect 259 478 361 524
use Inversor  Inversor_0 ~/icdesign/mag/Inversor
timestamp 1648588024
transform 1 0 335 0 1 478
box 0 0 608 984
use NAND  NAND_0 ~/icdesign/mag/NAND
timestamp 1648588519
transform 1 0 -327 0 1 478
box 0 0 608 984
use via  via_0 ~/icdesign/mag/Via
timestamp 1647641870
transform 1 0 398 0 1 712
box 31 179 97 245
<< end >>
